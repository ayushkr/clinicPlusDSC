




<svg height="210" width="500">
            <polygon points="200,10 250,190 160,{{:id}}" style="fill:lime;stroke:purple;stroke-width:1" />
            Sorry, your browser does not support inline SVG.

            <text x="0" y="15" fill="red">I love SVG!</text>
          </svg>

id={{:id}}


